package virtual_interface;
//    typedef virtual fifo_ifc.TB_Fifo vFIFO_T;
    typedef virtual cpu_ifc.TB_Sys2Dec vCPU_T;
    typedef virtual dec_ifc.TB_Dec2Bnc vDEC_T;
endpackage:virtual_interface
    
